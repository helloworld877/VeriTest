module and19 (
    input wire a,
    output wire out
);

assign out = &a;

endmodule
