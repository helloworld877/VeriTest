module decoder27 (d_out, d_in);

    output [15:0] d_out;
    input [3:0]   d_in;

assign d_out = (d_in == 4'b0000) ? (16'b0000_0000_0000_0001):
            (d_in == 4'b0001) ? (16'b0000_0000_0000_0001<<1):
            (d_in == 4'b0010) ? (16'b0000_0000_0000_0001<<2):
            (d_in == 4'b0011) ? (16'b0000_0000_0000_0001<<3):
            (d_in == 4'b0100) ? (16'b0000_0000_0000_0001<<4):
            (d_in == 4'b0101) ? (16'b0000_0000_0000_0001<<5):
            (d_in == 4'b0110) ? (16'b0000_0000_0000_0001<<6):
            (d_in == 4'b0111) ? (16'b0000_0000_0000_0001<<7):
            (d_in == 4'b1000) ? (16'b0000_0000_0000_0001<<8):
            (d_in == 4'b1001) ? (16'b0000_0000_0000_0001<<9):
            (d_in == 4'b1010) ? (16'b0000_0000_0000_0001<<10):
            (d_in == 4'b1011) ? (16'b0000_0000_0000_0001<<11):
            (d_in == 4'b1100) ? (16'b0000_0000_0000_0001<<12):
            (d_in == 4'b1101) ? (16'b0000_0000_0000_0001<<13):
            (d_in == 4'b1110) ? (16'b0000_0000_0000_0001<<14):
            (d_in == 4'b1111) ? (16'b0000_0000_0000_0001<<15):
	        16'b0000_0000_0000_0000;

endmodule