
module model(
    input A,
    input B,
    input C,
    output OUT
);
always @(*) begin
    
end
assign OUT = A&B&C;

endmodule
