module and_test (
    input wire a,
    output wire out
);

assign out = &a;

endmodule
