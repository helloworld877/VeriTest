//built-in operator
module or1 (
  input a,
  input b,
  output out
);

  assign out = a | b;

endmodule