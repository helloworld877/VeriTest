module not1 (
  input in,
  output out
);

  assign out = ~in; // Invert the input

endmodule