module or_gate(
  in4,in6, out
);


input in4, in6;
output out;

always @(*) begin
  
end
assign out = in4 | in6;

endmodule
