module not2 (
  input in,
  output out
);

  not (out, in); // Instantiate a NOT gate primitive

endmodule